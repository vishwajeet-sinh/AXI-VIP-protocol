class axi_sqr extends uvm_sequencer#(axi_tx);
    `uvm_component_utils(axi_sqr)
    `NEW
endclass